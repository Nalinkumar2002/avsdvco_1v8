magic
tech sky130A
timestamp 1628854847
<< nwell >>
rect -156 55 1139 56
rect -266 -373 1139 55
rect -266 -374 249 -373
rect -266 -376 -28 -374
<< nmos >>
rect 32 -505 50 -455
rect 168 -505 186 -455
rect 304 -504 322 -454
rect 440 -504 458 -454
rect 576 -504 594 -454
rect -133 -713 -115 -612
rect 784 -597 802 -453
rect 923 -518 941 -453
rect 32 -742 50 -613
rect 168 -742 186 -613
rect 304 -742 322 -613
rect 440 -742 458 -613
rect 576 -742 594 -613
<< pmos >>
rect -134 -190 -116 -89
rect 33 -190 51 -60
rect 169 -190 187 -60
rect 305 -190 323 -60
rect 441 -190 459 -60
rect 577 -190 595 -60
rect 32 -347 50 -297
rect 168 -347 186 -297
rect 304 -346 322 -296
rect 440 -346 458 -296
rect 576 -346 594 -296
rect 784 -346 802 -58
rect 923 -346 941 -217
<< ndiff >>
rect -13 -471 32 -455
rect -13 -489 -4 -471
rect 14 -489 32 -471
rect -13 -505 32 -489
rect 50 -471 95 -455
rect 50 -489 68 -471
rect 86 -489 95 -471
rect 50 -505 95 -489
rect 123 -471 168 -455
rect 123 -489 132 -471
rect 150 -489 168 -471
rect 123 -505 168 -489
rect 186 -471 231 -455
rect 186 -489 204 -471
rect 222 -489 231 -471
rect 186 -505 231 -489
rect 259 -470 304 -454
rect 259 -488 268 -470
rect 286 -488 304 -470
rect 259 -504 304 -488
rect 322 -470 367 -454
rect 322 -488 340 -470
rect 358 -488 367 -470
rect 322 -504 367 -488
rect 395 -470 440 -454
rect 395 -488 404 -470
rect 422 -488 440 -470
rect 395 -504 440 -488
rect 458 -470 503 -454
rect 458 -488 476 -470
rect 494 -488 503 -470
rect 458 -504 503 -488
rect 531 -470 576 -454
rect 531 -488 540 -470
rect 558 -488 576 -470
rect 531 -504 576 -488
rect 594 -470 639 -454
rect 594 -488 612 -470
rect 630 -488 639 -470
rect 594 -504 639 -488
rect 739 -462 784 -453
rect 739 -480 748 -462
rect 766 -480 784 -462
rect 739 -497 784 -480
rect 739 -514 748 -497
rect 766 -514 784 -497
rect 739 -531 784 -514
rect 739 -548 748 -531
rect 766 -548 784 -531
rect 739 -568 784 -548
rect 739 -585 748 -568
rect 766 -585 784 -568
rect -178 -632 -133 -612
rect -178 -650 -169 -632
rect -151 -650 -133 -632
rect -178 -673 -133 -650
rect -178 -691 -169 -673
rect -151 -691 -133 -673
rect -178 -713 -133 -691
rect -115 -633 -70 -612
rect 739 -597 784 -585
rect 802 -461 847 -453
rect 802 -479 820 -461
rect 838 -479 847 -461
rect 802 -497 847 -479
rect 802 -514 820 -497
rect 838 -514 847 -497
rect 802 -531 847 -514
rect 878 -470 923 -453
rect 878 -488 887 -470
rect 905 -488 923 -470
rect 878 -518 923 -488
rect 941 -470 986 -453
rect 941 -488 959 -470
rect 977 -488 986 -470
rect 941 -518 986 -488
rect 802 -548 820 -531
rect 838 -548 847 -531
rect 802 -568 847 -548
rect 802 -585 820 -568
rect 838 -585 847 -568
rect 802 -597 847 -585
rect -115 -650 -97 -633
rect -79 -650 -70 -633
rect -115 -675 -70 -650
rect -115 -692 -97 -675
rect -79 -692 -70 -675
rect -115 -713 -70 -692
rect -13 -633 32 -613
rect -13 -650 -3 -633
rect 15 -650 32 -633
rect -13 -671 32 -650
rect -13 -689 -4 -671
rect 14 -689 32 -671
rect -13 -709 32 -689
rect -13 -727 -4 -709
rect 14 -727 32 -709
rect -13 -742 32 -727
rect 50 -633 95 -613
rect 50 -650 68 -633
rect 86 -650 95 -633
rect 50 -673 95 -650
rect 50 -690 68 -673
rect 86 -690 95 -673
rect 50 -710 95 -690
rect 50 -727 68 -710
rect 86 -727 95 -710
rect 50 -742 95 -727
rect 123 -633 168 -613
rect 123 -650 133 -633
rect 151 -650 168 -633
rect 123 -671 168 -650
rect 123 -689 132 -671
rect 150 -689 168 -671
rect 123 -709 168 -689
rect 123 -727 132 -709
rect 150 -727 168 -709
rect 123 -742 168 -727
rect 186 -633 231 -613
rect 186 -650 204 -633
rect 222 -650 231 -633
rect 186 -673 231 -650
rect 186 -690 204 -673
rect 222 -690 231 -673
rect 186 -710 231 -690
rect 186 -727 204 -710
rect 222 -727 231 -710
rect 186 -742 231 -727
rect 259 -633 304 -613
rect 259 -650 269 -633
rect 287 -650 304 -633
rect 259 -671 304 -650
rect 259 -689 268 -671
rect 286 -689 304 -671
rect 259 -709 304 -689
rect 259 -727 268 -709
rect 286 -727 304 -709
rect 259 -742 304 -727
rect 322 -633 367 -613
rect 322 -650 340 -633
rect 358 -650 367 -633
rect 322 -673 367 -650
rect 322 -690 340 -673
rect 358 -690 367 -673
rect 322 -710 367 -690
rect 322 -727 340 -710
rect 358 -727 367 -710
rect 322 -742 367 -727
rect 395 -633 440 -613
rect 395 -650 405 -633
rect 423 -650 440 -633
rect 395 -671 440 -650
rect 395 -689 404 -671
rect 422 -689 440 -671
rect 395 -709 440 -689
rect 395 -727 404 -709
rect 422 -727 440 -709
rect 395 -742 440 -727
rect 458 -633 503 -613
rect 458 -650 476 -633
rect 494 -650 503 -633
rect 458 -673 503 -650
rect 458 -690 476 -673
rect 494 -690 503 -673
rect 458 -710 503 -690
rect 458 -727 476 -710
rect 494 -727 503 -710
rect 458 -742 503 -727
rect 531 -633 576 -613
rect 531 -650 541 -633
rect 559 -650 576 -633
rect 531 -671 576 -650
rect 531 -689 540 -671
rect 558 -689 576 -671
rect 531 -709 576 -689
rect 531 -727 540 -709
rect 558 -727 576 -709
rect 531 -742 576 -727
rect 594 -633 639 -613
rect 594 -650 612 -633
rect 630 -650 639 -633
rect 594 -673 639 -650
rect 594 -690 612 -673
rect 630 -690 639 -673
rect 594 -710 639 -690
rect 594 -727 612 -710
rect 630 -727 639 -710
rect 594 -742 639 -727
<< pdiff >>
rect -12 -75 33 -60
rect -179 -110 -134 -89
rect -179 -128 -170 -110
rect -152 -128 -134 -110
rect -179 -151 -134 -128
rect -179 -169 -170 -151
rect -152 -169 -134 -151
rect -179 -190 -134 -169
rect -116 -121 -71 -89
rect -116 -139 -97 -121
rect -79 -139 -71 -121
rect -116 -156 -71 -139
rect -116 -174 -98 -156
rect -80 -174 -71 -156
rect -116 -190 -71 -174
rect -12 -93 -3 -75
rect 15 -93 33 -75
rect -12 -113 33 -93
rect -12 -131 -3 -113
rect 15 -131 33 -113
rect -12 -152 33 -131
rect -12 -169 -2 -152
rect 16 -169 33 -152
rect -12 -190 33 -169
rect 51 -75 96 -60
rect 51 -92 69 -75
rect 87 -92 96 -75
rect 51 -112 96 -92
rect 51 -129 69 -112
rect 87 -129 96 -112
rect 51 -152 96 -129
rect 51 -169 69 -152
rect 87 -169 96 -152
rect 51 -190 96 -169
rect 124 -75 169 -60
rect 124 -93 133 -75
rect 151 -93 169 -75
rect 124 -113 169 -93
rect 124 -131 133 -113
rect 151 -131 169 -113
rect 124 -152 169 -131
rect 124 -169 134 -152
rect 152 -169 169 -152
rect 124 -190 169 -169
rect 187 -75 232 -60
rect 187 -92 205 -75
rect 223 -92 232 -75
rect 187 -112 232 -92
rect 187 -129 205 -112
rect 223 -129 232 -112
rect 187 -152 232 -129
rect 187 -169 205 -152
rect 223 -169 232 -152
rect 187 -190 232 -169
rect 260 -75 305 -60
rect 260 -93 269 -75
rect 287 -93 305 -75
rect 260 -113 305 -93
rect 260 -131 269 -113
rect 287 -131 305 -113
rect 260 -152 305 -131
rect 260 -169 270 -152
rect 288 -169 305 -152
rect 260 -190 305 -169
rect 323 -75 368 -60
rect 323 -92 341 -75
rect 359 -92 368 -75
rect 323 -112 368 -92
rect 323 -129 341 -112
rect 359 -129 368 -112
rect 323 -152 368 -129
rect 323 -169 341 -152
rect 359 -169 368 -152
rect 323 -190 368 -169
rect 396 -75 441 -60
rect 396 -93 405 -75
rect 423 -93 441 -75
rect 396 -113 441 -93
rect 396 -131 405 -113
rect 423 -131 441 -113
rect 396 -152 441 -131
rect 396 -169 406 -152
rect 424 -169 441 -152
rect 396 -190 441 -169
rect 459 -75 504 -60
rect 459 -92 477 -75
rect 495 -92 504 -75
rect 459 -112 504 -92
rect 459 -129 477 -112
rect 495 -129 504 -112
rect 459 -152 504 -129
rect 459 -169 477 -152
rect 495 -169 504 -152
rect 459 -190 504 -169
rect 532 -75 577 -60
rect 532 -93 541 -75
rect 559 -93 577 -75
rect 532 -113 577 -93
rect 532 -131 541 -113
rect 559 -131 577 -113
rect 532 -152 577 -131
rect 532 -169 542 -152
rect 560 -169 577 -152
rect 532 -190 577 -169
rect 595 -75 640 -60
rect 595 -92 613 -75
rect 631 -92 640 -75
rect 595 -112 640 -92
rect 595 -129 613 -112
rect 631 -129 640 -112
rect 595 -152 640 -129
rect 595 -169 613 -152
rect 631 -169 640 -152
rect 595 -190 640 -169
rect 739 -67 784 -58
rect 739 -85 748 -67
rect 766 -85 784 -67
rect 739 -102 784 -85
rect 739 -120 748 -102
rect 766 -120 784 -102
rect 739 -137 784 -120
rect 739 -155 748 -137
rect 766 -155 784 -137
rect 739 -172 784 -155
rect 739 -190 748 -172
rect 766 -190 784 -172
rect 739 -207 784 -190
rect 739 -225 748 -207
rect 766 -225 784 -207
rect 739 -242 784 -225
rect 739 -260 748 -242
rect 766 -260 784 -242
rect 739 -277 784 -260
rect 739 -295 748 -277
rect 766 -295 784 -277
rect -13 -313 32 -297
rect -13 -331 -4 -313
rect 14 -331 32 -313
rect -13 -347 32 -331
rect 50 -313 95 -297
rect 50 -331 68 -313
rect 86 -331 95 -313
rect 50 -347 95 -331
rect 123 -313 168 -297
rect 123 -331 132 -313
rect 150 -331 168 -313
rect 123 -347 168 -331
rect 186 -313 231 -297
rect 186 -331 204 -313
rect 222 -331 231 -313
rect 186 -347 231 -331
rect 259 -312 304 -296
rect 259 -330 268 -312
rect 286 -330 304 -312
rect 259 -346 304 -330
rect 322 -312 367 -296
rect 322 -330 340 -312
rect 358 -330 367 -312
rect 322 -346 367 -330
rect 395 -312 440 -296
rect 395 -330 404 -312
rect 422 -330 440 -312
rect 395 -346 440 -330
rect 458 -312 503 -296
rect 458 -330 476 -312
rect 494 -330 503 -312
rect 458 -346 503 -330
rect 531 -312 576 -296
rect 531 -330 540 -312
rect 558 -330 576 -312
rect 531 -346 576 -330
rect 594 -312 639 -296
rect 594 -330 612 -312
rect 630 -330 639 -312
rect 594 -346 639 -330
rect 739 -312 784 -295
rect 739 -330 748 -312
rect 766 -330 784 -312
rect 739 -346 784 -330
rect 802 -67 847 -58
rect 802 -85 821 -67
rect 839 -85 847 -67
rect 802 -102 847 -85
rect 802 -120 821 -102
rect 839 -120 847 -102
rect 802 -137 847 -120
rect 802 -155 821 -137
rect 839 -155 847 -137
rect 802 -172 847 -155
rect 802 -190 821 -172
rect 839 -190 847 -172
rect 802 -207 847 -190
rect 802 -225 821 -207
rect 839 -225 847 -207
rect 802 -242 847 -225
rect 802 -260 821 -242
rect 839 -260 847 -242
rect 802 -277 847 -260
rect 802 -295 821 -277
rect 839 -295 847 -277
rect 802 -312 847 -295
rect 802 -330 820 -312
rect 838 -330 847 -312
rect 802 -346 847 -330
rect 878 -242 923 -217
rect 878 -260 887 -242
rect 905 -260 923 -242
rect 878 -277 923 -260
rect 878 -295 887 -277
rect 905 -295 923 -277
rect 878 -312 923 -295
rect 878 -330 887 -312
rect 905 -330 923 -312
rect 878 -346 923 -330
rect 941 -241 986 -217
rect 941 -259 959 -241
rect 977 -259 986 -241
rect 941 -276 986 -259
rect 941 -294 959 -276
rect 977 -294 986 -276
rect 941 -312 986 -294
rect 941 -330 959 -312
rect 977 -330 986 -312
rect 941 -346 986 -330
<< ndiffc >>
rect -4 -489 14 -471
rect 68 -489 86 -471
rect 132 -489 150 -471
rect 204 -489 222 -471
rect 268 -488 286 -470
rect 340 -488 358 -470
rect 404 -488 422 -470
rect 476 -488 494 -470
rect 540 -488 558 -470
rect 612 -488 630 -470
rect 748 -480 766 -462
rect 748 -514 766 -497
rect 748 -548 766 -531
rect 748 -585 766 -568
rect -169 -650 -151 -632
rect -169 -691 -151 -673
rect 820 -479 838 -461
rect 820 -514 838 -497
rect 887 -488 905 -470
rect 959 -488 977 -470
rect 820 -548 838 -531
rect 820 -585 838 -568
rect -97 -650 -79 -633
rect -97 -692 -79 -675
rect -3 -650 15 -633
rect -4 -689 14 -671
rect -4 -727 14 -709
rect 68 -650 86 -633
rect 68 -690 86 -673
rect 68 -727 86 -710
rect 133 -650 151 -633
rect 132 -689 150 -671
rect 132 -727 150 -709
rect 204 -650 222 -633
rect 204 -690 222 -673
rect 204 -727 222 -710
rect 269 -650 287 -633
rect 268 -689 286 -671
rect 268 -727 286 -709
rect 340 -650 358 -633
rect 340 -690 358 -673
rect 340 -727 358 -710
rect 405 -650 423 -633
rect 404 -689 422 -671
rect 404 -727 422 -709
rect 476 -650 494 -633
rect 476 -690 494 -673
rect 476 -727 494 -710
rect 541 -650 559 -633
rect 540 -689 558 -671
rect 540 -727 558 -709
rect 612 -650 630 -633
rect 612 -690 630 -673
rect 612 -727 630 -710
<< pdiffc >>
rect -170 -128 -152 -110
rect -170 -169 -152 -151
rect -97 -139 -79 -121
rect -98 -174 -80 -156
rect -3 -93 15 -75
rect -3 -131 15 -113
rect -2 -169 16 -152
rect 69 -92 87 -75
rect 69 -129 87 -112
rect 69 -169 87 -152
rect 133 -93 151 -75
rect 133 -131 151 -113
rect 134 -169 152 -152
rect 205 -92 223 -75
rect 205 -129 223 -112
rect 205 -169 223 -152
rect 269 -93 287 -75
rect 269 -131 287 -113
rect 270 -169 288 -152
rect 341 -92 359 -75
rect 341 -129 359 -112
rect 341 -169 359 -152
rect 405 -93 423 -75
rect 405 -131 423 -113
rect 406 -169 424 -152
rect 477 -92 495 -75
rect 477 -129 495 -112
rect 477 -169 495 -152
rect 541 -93 559 -75
rect 541 -131 559 -113
rect 542 -169 560 -152
rect 613 -92 631 -75
rect 613 -129 631 -112
rect 613 -169 631 -152
rect 748 -85 766 -67
rect 748 -120 766 -102
rect 748 -155 766 -137
rect 748 -190 766 -172
rect 748 -225 766 -207
rect 748 -260 766 -242
rect 748 -295 766 -277
rect -4 -331 14 -313
rect 68 -331 86 -313
rect 132 -331 150 -313
rect 204 -331 222 -313
rect 268 -330 286 -312
rect 340 -330 358 -312
rect 404 -330 422 -312
rect 476 -330 494 -312
rect 540 -330 558 -312
rect 612 -330 630 -312
rect 748 -330 766 -312
rect 821 -85 839 -67
rect 821 -120 839 -102
rect 821 -155 839 -137
rect 821 -190 839 -172
rect 821 -225 839 -207
rect 821 -260 839 -242
rect 821 -295 839 -277
rect 820 -330 838 -312
rect 887 -260 905 -242
rect 887 -295 905 -277
rect 887 -330 905 -312
rect 959 -259 977 -241
rect 959 -294 977 -276
rect 959 -330 977 -312
<< psubdiff >>
rect -63 -812 -51 -794
rect -33 -812 -21 -794
rect 98 -812 110 -794
rect 128 -812 140 -794
rect 233 -812 245 -794
rect 263 -812 275 -794
rect 369 -812 381 -794
rect 399 -812 411 -794
rect 506 -812 518 -794
rect 536 -812 548 -794
rect 677 -812 689 -794
rect 707 -812 719 -794
rect 815 -812 827 -794
rect 845 -812 857 -794
<< nsubdiff >>
rect 121 10 170 12
rect -53 -8 -41 10
rect -23 -8 -11 10
rect 121 -8 135 10
rect 153 -8 170 10
rect 121 -13 170 -8
rect 261 -9 273 9
rect 291 -9 303 9
rect 390 -9 402 9
rect 420 -9 432 9
rect 525 -9 537 9
rect 555 -9 567 9
rect 679 -9 691 9
rect 709 -9 721 9
rect 808 -9 820 9
rect 838 -9 850 9
<< psubdiffcont >>
rect -51 -812 -33 -794
rect 110 -812 128 -794
rect 245 -812 263 -794
rect 381 -812 399 -794
rect 518 -812 536 -794
rect 689 -812 707 -794
rect 827 -812 845 -794
<< nsubdiffcont >>
rect -41 -8 -23 10
rect 135 -8 153 10
rect 273 -9 291 9
rect 402 -9 420 9
rect 537 -9 555 9
rect 691 -9 709 9
rect 820 -9 838 9
<< poly >>
rect 33 -60 51 -47
rect 169 -60 187 -47
rect 305 -60 323 -47
rect 441 -60 459 -47
rect 577 -60 595 -47
rect 784 -58 802 -45
rect -134 -89 -116 -76
rect -134 -206 -116 -190
rect 33 -206 51 -190
rect 169 -206 187 -190
rect 305 -206 323 -190
rect 441 -206 459 -190
rect 577 -206 595 -190
rect -134 -212 -98 -206
rect 33 -212 69 -206
rect 169 -212 205 -206
rect 305 -212 341 -206
rect 441 -212 477 -206
rect 577 -212 613 -206
rect -134 -214 -93 -212
rect -134 -232 -123 -214
rect -105 -232 -93 -214
rect -134 -234 -93 -232
rect 33 -214 74 -212
rect 33 -232 44 -214
rect 62 -232 74 -214
rect 33 -234 74 -232
rect 169 -214 210 -212
rect 169 -232 180 -214
rect 198 -232 210 -214
rect 169 -234 210 -232
rect 305 -214 346 -212
rect 305 -232 316 -214
rect 334 -232 346 -214
rect 305 -234 346 -232
rect 441 -214 482 -212
rect 441 -232 452 -214
rect 470 -232 482 -214
rect 441 -234 482 -232
rect 577 -214 618 -212
rect 577 -232 588 -214
rect 606 -232 618 -214
rect 577 -234 618 -232
rect -134 -240 -98 -234
rect 33 -240 69 -234
rect 169 -240 205 -234
rect 305 -240 341 -234
rect 441 -240 477 -234
rect 577 -240 613 -234
rect 32 -297 50 -279
rect 168 -297 186 -279
rect 304 -296 322 -278
rect 440 -296 458 -278
rect 576 -296 594 -278
rect 923 -217 941 -204
rect 32 -381 50 -347
rect 168 -381 186 -347
rect 304 -380 322 -346
rect 440 -380 458 -346
rect 576 -380 594 -346
rect 784 -380 802 -346
rect 923 -380 941 -346
rect 13 -387 50 -381
rect 149 -387 186 -381
rect 285 -386 322 -380
rect 421 -386 458 -380
rect 557 -386 594 -380
rect 765 -386 802 -380
rect 904 -386 941 -380
rect 8 -389 50 -387
rect 8 -407 20 -389
rect 38 -407 50 -389
rect 8 -409 50 -407
rect 144 -389 186 -387
rect 144 -407 156 -389
rect 174 -407 186 -389
rect 144 -409 186 -407
rect 280 -388 322 -386
rect 280 -406 292 -388
rect 310 -406 322 -388
rect 280 -408 322 -406
rect 416 -388 458 -386
rect 416 -406 428 -388
rect 446 -406 458 -388
rect 416 -408 458 -406
rect 552 -388 594 -386
rect 552 -406 564 -388
rect 582 -406 594 -388
rect 552 -408 594 -406
rect 760 -388 802 -386
rect 760 -406 772 -388
rect 790 -406 802 -388
rect 760 -408 802 -406
rect 899 -388 941 -386
rect 899 -406 911 -388
rect 929 -406 941 -388
rect 899 -408 941 -406
rect 13 -415 50 -409
rect 149 -415 186 -409
rect 285 -414 322 -408
rect 421 -414 458 -408
rect 557 -414 594 -408
rect 765 -414 802 -408
rect 904 -414 941 -408
rect 32 -455 50 -415
rect 168 -455 186 -415
rect 304 -454 322 -414
rect 440 -454 458 -414
rect 576 -454 594 -414
rect 784 -453 802 -414
rect 923 -453 941 -414
rect 32 -523 50 -505
rect 168 -523 186 -505
rect 304 -522 322 -504
rect 440 -522 458 -504
rect 576 -522 594 -504
rect -133 -568 -97 -562
rect 32 -568 68 -562
rect 168 -568 204 -562
rect 304 -568 340 -562
rect 440 -568 476 -562
rect 576 -568 612 -562
rect -133 -570 -92 -568
rect -133 -588 -122 -570
rect -104 -588 -92 -570
rect -133 -590 -92 -588
rect 32 -570 73 -568
rect 32 -588 43 -570
rect 61 -588 73 -570
rect 32 -590 73 -588
rect 168 -570 209 -568
rect 168 -588 179 -570
rect 197 -588 209 -570
rect 168 -590 209 -588
rect 304 -570 345 -568
rect 304 -588 315 -570
rect 333 -588 345 -570
rect 304 -590 345 -588
rect 440 -570 481 -568
rect 440 -588 451 -570
rect 469 -588 481 -570
rect 440 -590 481 -588
rect 576 -570 617 -568
rect 576 -588 587 -570
rect 605 -588 617 -570
rect 576 -590 617 -588
rect -133 -596 -97 -590
rect 32 -596 68 -590
rect 168 -596 204 -590
rect 304 -596 340 -590
rect 440 -596 476 -590
rect 576 -596 612 -590
rect -133 -612 -115 -596
rect 32 -613 50 -596
rect 168 -613 186 -596
rect 304 -613 322 -596
rect 440 -613 458 -596
rect 576 -613 594 -596
rect 923 -531 941 -518
rect 784 -610 802 -597
rect -133 -726 -115 -713
rect 32 -755 50 -742
rect 168 -755 186 -742
rect 304 -755 322 -742
rect 440 -755 458 -742
rect 576 -755 594 -742
<< polycont >>
rect -123 -232 -105 -214
rect 44 -232 62 -214
rect 180 -232 198 -214
rect 316 -232 334 -214
rect 452 -232 470 -214
rect 588 -232 606 -214
rect 20 -407 38 -389
rect 156 -407 174 -389
rect 292 -406 310 -388
rect 428 -406 446 -388
rect 564 -406 582 -388
rect 772 -406 790 -388
rect 911 -406 929 -388
rect -122 -588 -104 -570
rect 43 -588 61 -570
rect 179 -588 197 -570
rect 315 -588 333 -570
rect 451 -588 469 -570
rect 587 -588 605 -570
<< locali >>
rect -132 17 637 18
rect -132 10 920 17
rect -132 -8 -100 10
rect -82 -8 -41 10
rect -23 -8 70 10
rect 88 -8 135 10
rect 153 -8 206 10
rect 224 9 341 10
rect 224 -8 273 9
rect -132 -9 273 -8
rect 291 -8 341 9
rect 359 9 920 10
rect 359 -8 402 9
rect 291 -9 402 -8
rect 420 -9 477 9
rect 495 -9 537 9
rect 555 8 691 9
rect 555 -9 614 8
rect -132 -10 614 -9
rect 632 -9 691 8
rect 709 8 820 9
rect 709 -9 749 8
rect 632 -10 749 -9
rect 767 -9 820 8
rect 838 8 920 9
rect 838 -9 887 8
rect 767 -10 887 -9
rect 905 -10 920 8
rect -132 -19 920 -10
rect -178 -110 -144 -98
rect -178 -128 -170 -110
rect -152 -128 -144 -110
rect -178 -151 -144 -128
rect -178 -169 -170 -151
rect -152 -169 -144 -151
rect -178 -188 -144 -169
rect -106 -121 -74 -19
rect 61 -20 920 -19
rect 62 -60 96 -20
rect -106 -139 -97 -121
rect -79 -139 -74 -121
rect -106 -156 -74 -139
rect -106 -174 -98 -156
rect -80 -174 -74 -156
rect -106 -184 -74 -174
rect -11 -75 24 -60
rect -11 -93 -3 -75
rect 15 -93 24 -75
rect -11 -113 24 -93
rect -11 -131 -3 -113
rect 15 -131 24 -113
rect -11 -152 24 -131
rect -11 -169 -2 -152
rect 16 -169 24 -152
rect -178 -190 -146 -188
rect -11 -189 24 -169
rect 61 -75 95 -60
rect 61 -92 69 -75
rect 87 -92 95 -75
rect 61 -112 95 -92
rect 61 -129 69 -112
rect 87 -129 95 -112
rect 61 -152 95 -129
rect 61 -169 69 -152
rect 87 -169 95 -152
rect 61 -182 95 -169
rect 125 -75 160 -60
rect 125 -93 133 -75
rect 151 -93 160 -75
rect 125 -113 160 -93
rect 125 -131 133 -113
rect 151 -131 160 -113
rect 125 -152 160 -131
rect 125 -169 134 -152
rect 152 -169 160 -152
rect 125 -189 160 -169
rect 197 -75 231 -20
rect 197 -92 205 -75
rect 223 -92 231 -75
rect 197 -112 231 -92
rect 197 -129 205 -112
rect 223 -129 231 -112
rect 197 -152 231 -129
rect 197 -169 205 -152
rect 223 -169 231 -152
rect 197 -182 231 -169
rect 261 -75 296 -60
rect 261 -93 269 -75
rect 287 -93 296 -75
rect 261 -113 296 -93
rect 261 -131 269 -113
rect 287 -131 296 -113
rect 261 -152 296 -131
rect 261 -169 270 -152
rect 288 -169 296 -152
rect 261 -189 296 -169
rect 333 -75 367 -20
rect 470 -60 504 -20
rect 606 -60 640 -20
rect 333 -92 341 -75
rect 359 -92 367 -75
rect 333 -112 367 -92
rect 333 -129 341 -112
rect 359 -129 367 -112
rect 333 -152 367 -129
rect 333 -169 341 -152
rect 359 -169 367 -152
rect 333 -182 367 -169
rect 397 -75 432 -60
rect 397 -93 405 -75
rect 423 -93 432 -75
rect 397 -113 432 -93
rect 397 -131 405 -113
rect 423 -131 432 -113
rect 397 -152 432 -131
rect 397 -169 406 -152
rect 424 -169 432 -152
rect 397 -189 432 -169
rect 469 -61 504 -60
rect 469 -75 503 -61
rect 469 -92 477 -75
rect 495 -92 503 -75
rect 469 -112 503 -92
rect 469 -129 477 -112
rect 495 -129 503 -112
rect 469 -152 503 -129
rect 469 -169 477 -152
rect 495 -169 503 -152
rect 469 -182 503 -169
rect 533 -75 568 -60
rect 533 -93 541 -75
rect 559 -93 568 -75
rect 533 -113 568 -93
rect 533 -131 541 -113
rect 559 -131 568 -113
rect 533 -152 568 -131
rect 533 -169 542 -152
rect 560 -169 568 -152
rect 533 -189 568 -169
rect 605 -62 640 -60
rect 741 -62 775 -20
rect 605 -75 639 -62
rect 605 -92 613 -75
rect 631 -92 639 -75
rect 605 -112 639 -92
rect 605 -129 613 -112
rect 631 -129 639 -112
rect 605 -152 639 -129
rect 605 -169 613 -152
rect 631 -169 639 -152
rect 605 -182 639 -169
rect 740 -67 775 -62
rect 740 -85 748 -67
rect 766 -69 775 -67
rect 812 -67 844 -59
rect 766 -85 774 -69
rect 740 -102 774 -85
rect 740 -120 748 -102
rect 766 -120 774 -102
rect 740 -137 774 -120
rect 740 -155 748 -137
rect 766 -155 774 -137
rect 740 -172 774 -155
rect -175 -212 -146 -190
rect -6 -190 18 -189
rect 130 -190 154 -189
rect 266 -190 290 -189
rect 402 -190 426 -189
rect 538 -190 562 -189
rect 740 -190 748 -172
rect 766 -190 774 -172
rect -128 -212 -101 -206
rect -175 -214 -101 -212
rect -175 -232 -123 -214
rect -105 -232 -84 -214
rect -175 -237 -101 -232
rect -174 -622 -148 -237
rect -128 -240 -101 -237
rect -6 -305 17 -190
rect 39 -214 66 -206
rect 39 -232 44 -214
rect 62 -232 83 -214
rect 39 -240 66 -232
rect 130 -305 153 -190
rect 175 -214 202 -206
rect 175 -232 180 -214
rect 198 -232 219 -214
rect 175 -240 202 -232
rect 266 -304 289 -190
rect 311 -214 338 -206
rect 311 -232 316 -214
rect 334 -232 355 -214
rect 311 -240 338 -232
rect 402 -304 425 -190
rect 447 -214 474 -206
rect 447 -232 452 -214
rect 470 -232 491 -214
rect 447 -240 474 -232
rect 538 -304 561 -190
rect 583 -214 610 -206
rect 740 -207 774 -190
rect 583 -232 588 -214
rect 606 -232 627 -214
rect 740 -225 748 -207
rect 766 -225 774 -207
rect 583 -240 610 -232
rect 740 -242 774 -225
rect 740 -260 748 -242
rect 766 -260 774 -242
rect 740 -277 774 -260
rect 740 -295 748 -277
rect 766 -295 774 -277
rect -12 -313 22 -305
rect -12 -331 -4 -313
rect 14 -331 22 -313
rect -12 -341 22 -331
rect 60 -313 94 -306
rect 60 -331 68 -313
rect 86 -331 94 -313
rect 60 -347 94 -331
rect 124 -313 158 -305
rect 124 -331 132 -313
rect 150 -331 158 -313
rect 124 -341 158 -331
rect 196 -313 230 -306
rect 196 -331 204 -313
rect 222 -331 230 -313
rect 196 -347 230 -331
rect 260 -312 294 -304
rect 260 -330 268 -312
rect 286 -330 294 -312
rect 260 -340 294 -330
rect 332 -312 366 -305
rect 332 -330 340 -312
rect 358 -330 366 -312
rect 332 -346 366 -330
rect 396 -312 430 -304
rect 396 -330 404 -312
rect 422 -330 430 -312
rect 396 -340 430 -330
rect 468 -312 502 -305
rect 468 -330 476 -312
rect 494 -330 502 -312
rect 468 -346 502 -330
rect 532 -312 566 -304
rect 532 -330 540 -312
rect 558 -330 566 -312
rect 532 -340 566 -330
rect 604 -312 638 -305
rect 604 -330 612 -312
rect 630 -330 638 -312
rect 604 -346 638 -330
rect 740 -312 774 -295
rect 740 -330 748 -312
rect 766 -330 774 -312
rect 740 -340 774 -330
rect 812 -85 821 -67
rect 839 -85 844 -67
rect 812 -102 844 -85
rect 812 -120 821 -102
rect 839 -120 844 -102
rect 812 -137 844 -120
rect 812 -155 821 -137
rect 839 -155 844 -137
rect 812 -172 844 -155
rect 812 -190 821 -172
rect 839 -190 844 -172
rect 812 -207 844 -190
rect 812 -225 821 -207
rect 839 -225 844 -207
rect 812 -242 844 -225
rect 812 -260 821 -242
rect 839 -260 844 -242
rect 812 -277 844 -260
rect 812 -295 821 -277
rect 839 -295 844 -277
rect 812 -305 844 -295
rect 879 -242 913 -20
rect 879 -260 887 -242
rect 905 -260 913 -242
rect 879 -277 913 -260
rect 879 -295 887 -277
rect 905 -295 913 -277
rect 812 -312 846 -305
rect 812 -330 820 -312
rect 838 -330 846 -312
rect 812 -346 846 -330
rect 879 -312 913 -295
rect 879 -330 887 -312
rect 905 -330 913 -312
rect 879 -340 913 -330
rect 951 -241 985 -221
rect 951 -259 959 -241
rect 977 -259 985 -241
rect 951 -276 985 -259
rect 951 -294 959 -276
rect 977 -294 985 -276
rect 951 -312 985 -294
rect 951 -330 959 -312
rect 977 -330 985 -312
rect 951 -346 985 -330
rect 16 -389 43 -381
rect -1 -407 20 -389
rect 38 -407 43 -389
rect 16 -415 43 -407
rect 66 -389 88 -347
rect 152 -389 179 -381
rect 66 -407 156 -389
rect 174 -407 179 -389
rect 66 -455 88 -407
rect 152 -415 179 -407
rect 202 -389 224 -347
rect 288 -388 315 -380
rect 250 -389 292 -388
rect 202 -406 292 -389
rect 310 -406 315 -388
rect 202 -407 264 -406
rect 202 -455 224 -407
rect 288 -414 315 -406
rect 338 -388 360 -346
rect 424 -388 451 -380
rect 338 -406 428 -388
rect 446 -406 451 -388
rect 338 -454 360 -406
rect 424 -414 451 -406
rect 474 -388 496 -346
rect 560 -388 587 -380
rect 474 -406 564 -388
rect 582 -406 587 -388
rect 474 -454 496 -406
rect 560 -414 587 -406
rect 610 -388 632 -346
rect 768 -388 795 -380
rect 610 -406 645 -388
rect 666 -406 772 -388
rect 790 -406 795 -388
rect 610 -454 632 -406
rect 768 -414 795 -406
rect 818 -388 840 -346
rect 907 -388 934 -380
rect 818 -406 911 -388
rect 929 -406 934 -388
rect 818 -454 840 -406
rect 907 -414 934 -406
rect 957 -388 979 -346
rect 957 -406 999 -388
rect 957 -454 979 -406
rect -12 -471 22 -463
rect -12 -489 -4 -471
rect 14 -489 22 -471
rect -12 -499 22 -489
rect 60 -471 94 -455
rect 60 -489 68 -471
rect 86 -489 94 -471
rect 60 -497 94 -489
rect 124 -471 158 -463
rect 124 -489 132 -471
rect 150 -489 158 -471
rect 124 -499 158 -489
rect 196 -471 230 -455
rect 196 -489 204 -471
rect 222 -489 230 -471
rect 196 -497 230 -489
rect 260 -470 294 -462
rect 260 -488 268 -470
rect 286 -488 294 -470
rect 260 -498 294 -488
rect 332 -470 366 -454
rect 332 -488 340 -470
rect 358 -488 366 -470
rect 332 -496 366 -488
rect 396 -470 430 -462
rect 396 -488 404 -470
rect 422 -488 430 -470
rect 396 -498 430 -488
rect 468 -470 502 -454
rect 468 -488 476 -470
rect 494 -488 502 -470
rect 468 -496 502 -488
rect 532 -470 566 -462
rect 532 -488 540 -470
rect 558 -488 566 -470
rect 532 -498 566 -488
rect 604 -470 638 -454
rect 741 -462 774 -455
rect 604 -488 612 -470
rect 630 -488 638 -470
rect 604 -496 638 -488
rect 740 -480 748 -462
rect 766 -480 774 -462
rect 740 -497 774 -480
rect -127 -570 -100 -562
rect -127 -588 -122 -570
rect -104 -588 -83 -570
rect -127 -596 -100 -588
rect -7 -612 16 -499
rect 38 -570 65 -562
rect 38 -588 43 -570
rect 61 -588 82 -570
rect 38 -596 65 -588
rect 129 -612 152 -499
rect 174 -570 201 -562
rect 174 -588 179 -570
rect 197 -588 218 -570
rect 174 -596 201 -588
rect 265 -612 288 -498
rect 310 -570 337 -562
rect 310 -588 315 -570
rect 333 -588 354 -570
rect 310 -596 337 -588
rect 401 -612 424 -498
rect 446 -570 473 -562
rect 446 -588 451 -570
rect 469 -588 490 -570
rect 446 -596 473 -588
rect 537 -612 560 -498
rect 740 -514 748 -497
rect 766 -514 774 -497
rect 740 -531 774 -514
rect 740 -548 748 -531
rect 766 -548 774 -531
rect 582 -570 609 -562
rect 740 -568 774 -548
rect 582 -588 587 -570
rect 605 -588 626 -570
rect 740 -585 748 -568
rect 766 -585 774 -568
rect 812 -461 846 -454
rect 812 -479 820 -461
rect 838 -479 846 -461
rect 812 -497 846 -479
rect 812 -514 820 -497
rect 838 -514 846 -497
rect 879 -470 913 -462
rect 879 -488 887 -470
rect 905 -488 913 -470
rect 879 -498 913 -488
rect 951 -470 985 -454
rect 951 -488 959 -470
rect 977 -488 985 -470
rect 951 -496 985 -488
rect 812 -531 846 -514
rect 812 -548 820 -531
rect 838 -548 846 -531
rect 812 -568 846 -548
rect 812 -585 820 -568
rect 838 -585 846 -568
rect 582 -596 609 -588
rect -7 -613 17 -612
rect 129 -613 153 -612
rect 265 -613 289 -612
rect 401 -613 425 -612
rect 537 -613 561 -612
rect -177 -632 -142 -622
rect -177 -650 -169 -632
rect -151 -650 -142 -632
rect -177 -673 -142 -650
rect -177 -691 -169 -673
rect -151 -691 -142 -673
rect -177 -713 -142 -691
rect -105 -633 -71 -622
rect -105 -650 -97 -633
rect -79 -650 -71 -633
rect -105 -675 -71 -650
rect -105 -692 -97 -675
rect -79 -692 -71 -675
rect -105 -713 -71 -692
rect -12 -633 23 -613
rect -12 -650 -3 -633
rect 15 -650 23 -633
rect -12 -671 23 -650
rect -12 -689 -4 -671
rect 14 -689 23 -671
rect -12 -709 23 -689
rect -101 -784 -74 -713
rect -12 -727 -4 -709
rect 14 -727 23 -709
rect -12 -742 23 -727
rect 60 -633 94 -620
rect 60 -650 68 -633
rect 86 -650 94 -633
rect 60 -673 94 -650
rect 60 -690 68 -673
rect 86 -690 94 -673
rect 60 -710 94 -690
rect 60 -727 68 -710
rect 86 -727 94 -710
rect 60 -742 94 -727
rect 124 -633 159 -613
rect 124 -650 133 -633
rect 151 -650 159 -633
rect 124 -671 159 -650
rect 124 -689 132 -671
rect 150 -689 159 -671
rect 124 -709 159 -689
rect 124 -727 132 -709
rect 150 -727 159 -709
rect 124 -742 159 -727
rect 196 -633 230 -620
rect 196 -650 204 -633
rect 222 -650 230 -633
rect 196 -673 230 -650
rect 196 -690 204 -673
rect 222 -690 230 -673
rect 196 -710 230 -690
rect 196 -727 204 -710
rect 222 -727 230 -710
rect 196 -742 230 -727
rect 260 -633 295 -613
rect 260 -650 269 -633
rect 287 -650 295 -633
rect 260 -671 295 -650
rect 260 -689 268 -671
rect 286 -689 295 -671
rect 260 -709 295 -689
rect 260 -727 268 -709
rect 286 -727 295 -709
rect 260 -742 295 -727
rect 332 -633 366 -620
rect 332 -650 340 -633
rect 358 -650 366 -633
rect 332 -673 366 -650
rect 332 -690 340 -673
rect 358 -690 366 -673
rect 332 -710 366 -690
rect 332 -727 340 -710
rect 358 -727 366 -710
rect 332 -742 366 -727
rect 396 -633 431 -613
rect 396 -650 405 -633
rect 423 -650 431 -633
rect 396 -671 431 -650
rect 396 -689 404 -671
rect 422 -689 431 -671
rect 396 -709 431 -689
rect 396 -727 404 -709
rect 422 -727 431 -709
rect 396 -742 431 -727
rect 468 -633 502 -620
rect 468 -650 476 -633
rect 494 -650 502 -633
rect 468 -673 502 -650
rect 468 -690 476 -673
rect 494 -690 502 -673
rect 468 -710 502 -690
rect 468 -727 476 -710
rect 494 -727 502 -710
rect 468 -742 502 -727
rect 532 -633 567 -613
rect 532 -650 541 -633
rect 559 -650 567 -633
rect 532 -671 567 -650
rect 532 -689 540 -671
rect 558 -689 567 -671
rect 532 -709 567 -689
rect 532 -727 540 -709
rect 558 -727 567 -709
rect 532 -742 567 -727
rect 604 -633 638 -620
rect 604 -650 612 -633
rect 630 -650 638 -633
rect 604 -673 638 -650
rect 604 -690 612 -673
rect 630 -690 638 -673
rect 604 -710 638 -690
rect 604 -727 612 -710
rect 630 -727 638 -710
rect 604 -742 638 -727
rect 61 -784 93 -742
rect 197 -784 229 -742
rect 334 -784 366 -742
rect 469 -784 501 -742
rect 605 -784 637 -742
rect 740 -784 774 -585
rect 813 -589 846 -585
rect 881 -784 912 -498
rect -131 -794 934 -784
rect -131 -812 -98 -794
rect -80 -812 -51 -794
rect -33 -812 21 -794
rect 39 -812 110 -794
rect 128 -812 177 -794
rect 195 -812 245 -794
rect 263 -812 313 -794
rect 331 -812 381 -794
rect 399 -812 451 -794
rect 469 -812 518 -794
rect 536 -812 611 -794
rect 629 -812 689 -794
rect 707 -812 745 -794
rect 763 -812 827 -794
rect 845 -812 888 -794
rect 906 -812 934 -794
rect -131 -823 934 -812
<< viali >>
rect -100 -8 -82 10
rect 70 -8 88 10
rect 206 -8 224 10
rect 341 -8 359 10
rect 477 -9 495 9
rect 614 -10 632 8
rect 749 -10 767 8
rect 887 -10 905 8
rect -84 -232 -65 -214
rect 83 -232 102 -214
rect 219 -232 238 -214
rect 355 -232 374 -214
rect 491 -232 510 -214
rect 627 -232 646 -214
rect -22 -407 -1 -389
rect 645 -406 666 -388
rect 999 -406 1017 -388
rect -83 -588 -64 -570
rect 82 -588 101 -570
rect 218 -588 237 -570
rect 354 -588 373 -570
rect 490 -588 509 -570
rect 626 -588 645 -570
rect -98 -812 -80 -794
rect 21 -812 39 -794
rect 177 -812 195 -794
rect 313 -812 331 -794
rect 451 -812 469 -794
rect 611 -812 629 -794
rect 745 -812 763 -794
rect 888 -812 906 -794
<< metal1 >>
rect -132 10 919 18
rect -132 -8 -100 10
rect -82 -8 70 10
rect 88 -8 206 10
rect 224 -8 341 10
rect 359 9 919 10
rect 359 -8 477 9
rect -132 -9 477 -8
rect 495 8 919 9
rect 495 -9 614 8
rect -132 -10 614 -9
rect 632 -10 749 8
rect 767 -10 887 8
rect 905 -10 919 8
rect -132 -18 919 -10
rect -132 -19 58 -18
rect -134 -214 653 -209
rect -134 -232 -84 -214
rect -65 -232 83 -214
rect 102 -232 219 -214
rect 238 -232 355 -214
rect 374 -232 491 -214
rect 510 -232 627 -214
rect 646 -232 653 -214
rect -134 -238 653 -232
rect -28 -388 672 -383
rect -28 -389 645 -388
rect -28 -407 -22 -389
rect -1 -406 645 -389
rect 666 -406 672 -388
rect -1 -407 672 -406
rect -28 -412 672 -407
rect 984 -388 1040 -383
rect 984 -406 999 -388
rect 1017 -406 1040 -388
rect 984 -412 1040 -406
rect -133 -564 -97 -538
rect -133 -570 652 -564
rect -133 -588 -83 -570
rect -64 -588 82 -570
rect 101 -588 218 -570
rect 237 -588 354 -570
rect 373 -588 490 -570
rect 509 -588 626 -570
rect 645 -588 652 -570
rect -133 -593 652 -588
rect -132 -794 934 -783
rect -132 -812 -98 -794
rect -80 -812 21 -794
rect 39 -812 177 -794
rect 195 -812 313 -794
rect 331 -812 451 -794
rect 469 -812 611 -794
rect 629 -812 745 -794
rect 763 -812 888 -794
rect 906 -812 934 -794
rect -132 -824 934 -812
<< labels >>
flabel metal1 -126 -556 -104 -551 0 FreeSans 40 0 0 80 VCTRL
flabel metal1 -117 -10 -112 12 0 FreeSans 40 270 0 -80 VDD
flabel metal1 1021 -406 1024 -388 0 FreeSans 40 90 0 -80 F_OUT
flabel metal1 -114 -817 -109 -792 0 FreeSans 40 270 0 -80 GND
<< end >>
